module main();
    initial begin
        $display("Hello World");
    end
endmodule

